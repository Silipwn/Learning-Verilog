module fulladd(sum, c_out, a, b, c_in);

output[3:0] sum;
output c_cout;

input [3:0] a,b;

input c_in;

endmodule
