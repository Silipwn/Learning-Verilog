module Multi(x1,x2,c,f);
    input x1,x2,c;
    output f;

    not(k,s);
    and(g,k,x1);
    and(h,s,x2);
    or(f,g,h);
endmodule
