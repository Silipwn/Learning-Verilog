module adder(a,b,c,s);
    input a,b;
    output c,s;
    
    assign c = a&b;
    assign s = a^b;
endmodule

module sub(a,b,c,s);
    input(

module display(s0,s1,a,b,c,d,e,f,g);
    input s0,s1;
    output a,b,c,d,e,f,g;
    
